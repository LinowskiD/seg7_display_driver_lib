library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package defines_pkg is

  constant c_number_of_digits_default : natural := 4;

end package defines_pkg;